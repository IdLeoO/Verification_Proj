`ifndef DRIVER_SV
`define DRIVER_SV


class Driver;    
    

    
    extern function new(your code);
    extern task run();
    
    
endclass
 
function Driver::new(your code);
endfunction



task Driver::run();
endtask

`endif

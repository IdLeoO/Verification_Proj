`ifndef GEN_SV
`define GEN_SV


class Gen ;

extern function new(/*your code*/);
extern virtual task run();

endclass

function Gen::new(/*your code*/);
endfunction

task Gen::run();
endtask

`endif

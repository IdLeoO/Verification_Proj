`ifndef MONITOR_SV
`define MONITOR_SV


class Mon;
    
    extern function new(/*your code*/);
    extern task run();
endclass

function Mon::new(/*your code*/);
  
endfunction

task Mon::run();
    
endtask

`endif

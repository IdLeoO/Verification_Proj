`ifndef PACKAGE_SV
`define PACKAGE_SV

package chnl_pkg;





endpackage
`endif
 
`ifndef SCB_SV
`define SCB_SV

class Scb;
    
    extern function new(/*your code*/);
    extern task run();
endclass

function Scb::new(/*your code*/);

endfunction



task Scb::run();
            
endtask
`endif
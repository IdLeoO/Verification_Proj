module mcdf_property(
    // input interface
);

    //  Add assertion here

endmodule
`ifndef REF_MODEL_SV
`define REF_MODEL_SV


class Ref_model;    
    

    /*your code*/
    
    extern function new(/*your code*/);
    extern task run();


    
    
endclass
 
function Ref_model::new(/*your code*/);
   
endfunction

task Ref_model::run();

endtask



`endif


